library ieee;
use ieee.std_logic_1164.all;

--------------------------------------------------

entity k_reg is
port(k_out: out std_logic_vector (0 to 2047)
);
end k_reg;  

--------------------------------------------------

architecture k_reg_arch of k_reg is

begin
	k_out <= X"428A2F9871374491B5C0FBCFE9B5DBA53956C25B59F111F1923F82A4AB1C5ED5D807AA9812835B01243185BE550C7DC372BE5D7480DEB1FE9BDC06A7C19BF174E49B69C1EFBE47860FC19DC6240CA1CC2DE92C6F4A7484AA5CB0A9DC76F988DA983E5152A831C66DB00327C8BF597FC7C6E00BF3D5A7914706CA63511429296727B70A852E1B21384D2C6DFC53380D13650A7354766A0ABB81C2C92E92722C85A2BFE8A1A81A664BC24B8B70C76C51A3D192E819D6990624F40E3585106AA07019A4C1161E376C082748774C34B0BCB5391C0CB34ED8AA4A5B9CCA4F682E6FF3748F82EE78A5636F84C878148CC7020890BEFFFAA4506CEBBEF9A3F7C67178F2";
end k_reg_arch;